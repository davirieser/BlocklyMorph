$ 3 0.000005 382.76258214399064 50 5 50 5e-11
w 384 208 400 208 0
207 512 144 592 144 4 out
R 80 48 80 0 0 0 40 5 0 0 0.5
g 80 272 80 304 0 0
r 80 160 80 272 0 120000
w 64 144 80 144 0
r 80 48 80 144 0 330000
r 112 48 192 48 0 330000
r 192 112 192 176 0 120000
r 192 224 192 288 0 100000
g 192 288 192 304 0 0
w 80 48 112 48 0
w 192 176 192 192 0
w 192 192 192 224 0
w 192 224 224 224 0
w 176 192 224 192 0
a 256 96 368 96 9 5 0 1000000 1.3333333333333333 1.999999999986457 100000
w 192 80 256 80 0
w 192 112 192 80 0
w 192 80 192 48 0
w 176 112 256 112 0
a 256 208 368 208 9 5 0 1000000 0.9090909090847531 1.3333333333333333 100000
w 224 192 256 192 0
w 224 224 256 224 0
w 368 208 384 208 0
w 368 96 384 96 0
207 64 144 0 144 4 in
w 80 144 80 160 0
151 400 144 512 144 0 2 0 5
w 384 96 400 96 0
w 400 96 400 128 0
w 400 160 400 208 0
w 176 112 144 112 0
w 144 112 144 192 0
w 144 192 176 192 0
w 80 144 144 144 0
w 144 144 144 112 0
x 256 73 280 76 4 20 2V
x 238 246 279 249 4 20 0.9V
