$ 17 0.000005 382.76258214399064 50 5 50 5e-11
L 192 400 128 400 0 0 false 5 0
L 192 432 128 432 0 0 false 5 0
185 192 224 304 224 0 2
R 192 224 144 224 0 0 40 5 0 0 0.5
w 192 400 224 400 0
w 224 384 224 400 0
w 192 432 256 432 0
w 256 432 256 384 0
L 80 0 -48 0 0 1 false 5 0
. Window\sComparator 0 2 1 2 in 8 0 2 out 6 0 3 TransistorElm\s1\s2\s3\rTransistorElm\s4\s3\s0\rRailElm\s7\rResistorElm\s8\s0\rResistorElm\s7\s8\rResistorElm\s7\s9\rResistorElm\s9\s10\rResistorElm\s10\s0\rResistorElm\s11\s1\rResistorElm\s5\s4\rOpAmpElm\s8\s9\s11\rOpAmpElm\s10\s8\s5\rResistorElm\s2\s12\rRailElm\s12\rRailElm\s13\rResistorElm\s13\s6\rTransistorElm\s2\s6\s0 0\\s1\\s0.5700403623732102\\s0.6401396095088427\\s100\\sdefault\s0\\s1\\s0.5702234559618686\\s0.6420695171207146\\s100\\sdefault\s0\\s0\\s40\\s5\\s0\\s0\\s0.5\s0\\s120000\s0\\s330000\s0\\s330000\s0\\s120000\s0\\s100000\s0\\s10000\s0\\s10000\s9\\s5\\s0\\s1000000\\s1.3333333333333333\\s1.999999999986457\\s100000\s9\\s5\\s0\\s1000000\\s0.9090909090847531\\s1.3333333333333333\\s100000\s0\\s1000\s0\\s0\\s40\\s5\\s0\\s0\\s0.5\s0\\s0\\s40\\s5\\s0\\s0\\s0.5\s0\\s1000\s0\\s1\\s-4.8580546575718415\\s0.1419453082944785\\s100\\sdefault
410 256 0 400 0 1 Window\sComparator 0\s1\s-0.6629458831519461\s-0.018228241723234777\s100\sdefault 0\s1\s0.5738673613748971\s0.5917956132344714\s100\sdefault 0\s0\s40\s5\s0\s0\s0.5 0\s120000 0\s330000 0\s330000 0\s120000 0\s100000 0\s10000 0\s10000 9\s5\s0\s1000000\s5\s2.0000000000015112\s100000 9\s5\s0\s1000000\s0.909090909093635\s5\s100000 0\s1000 0\s0\s40\s5\s0\s0\s0.5 0\s0\s40\s5\s0\s0\s0.5 0\s1000 0\s1\s0.63270414458758\s0.6626458932882856\s100\sdefault
w 80 0 256 0 0
w 352 0 496 0 0
w 320 224 416 224 0
w 416 224 416 64 0
w 416 64 464 64 0
t 560 -16 560 -48 0 1 0 0 100 default
w 576 -48 592 -48 0
w 464 64 464 -16 0
w 544 -48 176 -48 0
w 176 -48 -32 -48 0
w 192 32 512 32 0
w 608 80 704 80 0
r 464 -16 560 -16 0 100000
r 592 -48 672 -48 0 1000
L 672 -48 720 -48 0 1 false 5 0
w 496 0 704 0 0
w 464 64 480 64 0
w 80 0 80 32 0
w 512 32 608 32 0
w 608 32 608 48 0
r 176 -48 176 -112 0 1000000
R 176 -112 176 -144 0 0 40 5 0 0 0.5
R 224 512 224 480 0 0 40 5 0 0 0.5
r 224 576 224 512 0 1000000
w 656 656 656 672 0
w 560 656 656 656 0
w 128 624 128 656 0
w 544 624 752 624 0
L 720 576 768 576 0 0 false 5 0
r 640 576 720 576 0 1000
r 512 608 608 608 0 100000
w 656 704 752 704 0
w 240 656 560 656 0
w 224 576 16 576 0
w 592 576 224 576 0
w 512 688 512 608 0
w 624 576 640 576 0
t 608 608 608 576 0 1 8.106370003019671e-23 -4.999994843905212 100 default
w 464 688 512 688 0
w 400 624 544 624 0
w 128 624 304 624 0
410 304 624 448 624 1 Window\sComparator 0\s1\s0.570040362373211\s0.6401396095088427\s100\sdefault 0\s1\s0.5702234559618673\s0.6420695171207146\s100\sdefault 0\s0\s40\s5\s0\s0\s0.5 0\s120000 0\s330000 0\s330000 0\s120000 0\s100000 0\s10000 0\s10000 9\s5\s0\s1000000\s1.3333333333331865\s1.9999999999686935\s100000 9\s5\s0\s1000000\s0.9090909090820884\s1.3333333333331865\s100000 0\s1000 0\s0\s40\s5\s0\s0\s0.5 0\s0\s40\s5\s0\s0\s0.5 0\s1000 0\s1\s-4.858054657571842\s0.14194530829447902\s100\sdefault
w 464 688 464 256 0
w 320 256 464 256 0
w 128 624 16 624 0
w 80 32 192 32 0
f 560 64 608 64 32 1.5 0.02
w 480 64 560 64 0
w 128 656 240 656 0
f 592 688 656 688 32 1.5 0.02
w 512 688 592 688 0

