$ 17 0.000005 382.76258214399064 50 5 50 5e-11
L 192 400 128 400 0 0 false 5 0
L 192 432 128 432 0 0 false 5 0
185 192 224 304 224 0 2
R 192 224 144 224 0 0 40 5 0 0 0.5
w 192 400 224 400 0
w 224 384 224 400 0
w 192 432 256 432 0
w 256 432 256 384 0
L 80 0 -48 0 0 1 false 5 0
. Window\sComparator 0 2 1 2 in 8 0 2 out 6 0 3 TransistorElm\s1\s2\s3\rTransistorElm\s4\s3\s0\rRailElm\s7\rResistorElm\s8\s0\rResistorElm\s7\s8\rResistorElm\s7\s9\rResistorElm\s9\s10\rResistorElm\s10\s0\rResistorElm\s11\s1\rResistorElm\s5\s4\rOpAmpElm\s8\s9\s11\rOpAmpElm\s10\s8\s5\rResistorElm\s2\s12\rRailElm\s12\rRailElm\s13\rResistorElm\s13\s6\rTransistorElm\s2\s6\s0 0\\s1\\s0.5700403623732102\\s0.6401396095088427\\s100\\sdefault\s0\\s1\\s0.5702234559618686\\s0.6420695171207146\\s100\\sdefault\s0\\s0\\s40\\s5\\s0\\s0\\s0.5\s0\\s120000\s0\\s330000\s0\\s330000\s0\\s120000\s0\\s100000\s0\\s10000\s0\\s10000\s9\\s5\\s0\\s1000000\\s1.3333333333333333\\s1.999999999986457\\s100000\s9\\s5\\s0\\s1000000\\s0.9090909090847531\\s1.3333333333333333\\s100000\s0\\s1000\s0\\s0\\s40\\s5\\s0\\s0\\s0.5\s0\\s0\\s40\\s5\\s0\\s0\\s0.5\s0\\s1000\s0\\s1\\s-4.8580546575718415\\s0.1419453082944785\\s100\\sdefault
410 256 0 400 0 1 Window\sComparator 0\s1\s-0.6629458831519461\s-0.018228241723234898\s100\sdefault 0\s1\s0.573867361374897\s0\s100\sdefault 0\s0\s40\s5\s0\s0\s0.5 0\s120000 0\s330000 0\s330000 0\s120000 0\s100000 0\s10000 0\s10000 9\s5\s0\s1000000\s5\s2.0000000000015112\s100000 9\s5\s0\s1000000\s0.909090909093635\s5\s100000 0\s1000 0\s0\s40\s5\s0\s0\s0.5 0\s0\s40\s5\s0\s0\s0.5 0\s1000 0\s1\s0.63270414458758\s0\s100\sdefault
w 80 0 256 0 0
w 352 0 496 0 0
w 320 224 416 224 0
w 416 224 416 64 0
w 416 -16 464 -16 0
t 560 -16 560 -48 0 1 0.5147567164084298 0.5114121891986025 100 default
w 576 -48 592 -48 0
w 416 64 416 -16 0
w 544 -48 176 -48 0
w 176 -48 -32 -48 0
r 464 -16 560 -16 0 100000
r 592 -48 672 -48 0 1000
L 672 -48 720 -48 0 1 false 5 0
w 496 0 704 0 0
w 80 0 80 32 0
r 176 -48 176 -112 0 1000000
R 176 -112 176 -144 0 0 40 5 0 0 0.5
R 224 512 224 480 0 0 40 5 0 0 0.5
r 224 576 224 512 0 1000000
w 128 624 128 656 0
w 544 624 752 624 0
L 720 576 768 576 0 0 false 5 0
r 640 576 720 576 0 1000
r 512 608 608 608 0 100000
w 224 576 16 576 0
w 592 576 224 576 0
w 624 576 640 576 0
t 608 608 608 576 0 1 0.009045039526561065 -4.990949762511912 100 default
w 400 624 544 624 0
410 304 624 448 624 1 Window\sComparator 0\s1\s0.5700403623732121\s0.6401396095088427\s100\sdefault 0\s1\s0.5702234559618645\s0\s100\sdefault 0\s0\s40\s5\s0\s0\s0.5 0\s120000 0\s330000 0\s330000 0\s120000 0\s100000 0\s10000 0\s10000 9\s5\s0\s1000000\s1.3333333333333333\s1.9999999999953388\s100000 9\s5\s0\s1000000\s0.9090909090847532\s1.3333333333333333\s100000 0\s1000 0\s0\s40\s5\s0\s0\s0.5 0\s0\s40\s5\s0\s0\s0.5 0\s1000 0\s1\s-4.858054657571841\s0\s100\sdefault
w 320 256 464 256 0
w 128 624 -48 624 0
w 80 32 192 32 0
w 128 656 240 656 0
184 864 240 1008 240 0 2
w 192 32 832 32 0
w 832 32 832 240 0
w 832 240 864 240 0
w 224 400 928 400 0
w 256 432 960 432 0
w 960 432 960 400 0
w 752 624 832 624 0
w 832 272 864 272 0
w 992 240 1152 240 0
w 128 624 304 624 0
w 240 656 816 656 0
w 816 656 816 272 0
w 816 272 832 272 0
x 756 -47 786 -44 4 24 TX
x 754 4 787 7 4 24 RX
x 863 631 896 634 4 24 RX
x 749 556 779 559 4 24 TX
x -131 4 -101 7 4 24 TX
x -126 -42 -93 -39 4 24 RX
x -69 580 -36 583 4 24 RX
x -119 628 -89 631 4 24 TX
