$ 17 0.000005 382.76258214399064 50 5 50 5e-11
t 496 96 528 96 0 1 0.5700403623732129 0.640139609508843 100 default
t 496 208 528 208 0 1 0.5702234559618667 0.6420695171207146 100 default
w 384 208 400 208 0
w 528 112 528 192 0
g 528 336 528 368 0 0
207 672 80 752 80 4 out
R 80 48 80 0 0 0 40 5 0 0 0.5
g 80 256 80 288 0 0
r 80 144 80 256 0 120000
w 64 144 80 144 0
w 80 144 176 144 0
w 176 144 176 112 0
r 80 48 80 144 0 330000
r 112 48 192 48 0 330000
r 192 112 192 176 0 120000
r 192 224 192 288 0 100000
g 192 288 192 304 0 0
w 80 48 112 48 0
w 192 176 192 192 0
w 192 192 192 224 0
r 384 96 480 96 0 10000
r 400 208 496 208 0 10000
w 528 224 528 256 0
w 192 224 224 224 0
w 176 144 176 192 0
w 176 192 224 192 0
a 256 96 368 96 9 5 0 1000000 1.3333333333333333 1.999999999986457 100000
w 192 80 256 80 0
w 192 112 192 80 0
w 192 80 192 48 0
w 176 112 256 112 0
a 256 208 368 208 9 5 0 1000000 0.9090909090847531 1.3333333333333333 100000
w 224 192 256 192 0
w 224 224 256 224 0
w 368 208 384 208 0
w 64 144 -32 144 0
w 368 96 384 96 0
w 480 96 496 96 0
w 528 256 528 336 0
r 528 80 528 0 0 1000
R 528 0 528 -48 0 0 40 5 0 0 0.5
R 592 0 592 -48 0 0 40 5 0 0 0.5
r 592 0 592 80 0 1000
t 560 96 592 96 0 1 -4.858054657571842 0.1419453082944779 100 default
w 528 80 560 80 0
w 560 80 560 96 0
w 528 256 592 256 0
w 592 112 592 256 0
w 592 80 672 80 0
207 -32 144 -96 144 4 in

